magic
tech sky130A
timestamp 1723068911
<< metal1 >>
rect 100 21000 9900 21200
rect 100 20840 300 21000
rect 100 20830 640 20840
rect 100 20780 240 20830
rect 290 20820 640 20830
rect 3260 20820 3680 20840
rect 290 20780 300 20820
rect 100 20700 300 20780
rect 3340 20790 3390 20800
rect 3340 20760 3350 20790
rect 3380 20780 3390 20790
rect 3380 20760 3600 20780
rect 4090 20770 4160 20780
rect 3340 20750 3390 20760
rect 4090 20730 4100 20770
rect 4010 20720 4100 20730
rect 4150 20720 4160 20770
rect 4010 20710 4160 20720
rect 4190 20770 4260 20780
rect 4190 20720 4200 20770
rect 4250 20720 4260 20770
rect 4190 20710 4260 20720
rect 3940 20660 4410 20680
rect 230 18230 640 18240
rect 230 18180 240 18230
rect 290 18220 640 18230
rect 3260 18220 3690 18240
rect 290 18180 300 18220
rect 230 18170 300 18180
rect 3340 18190 3390 18200
rect 3340 18160 3350 18190
rect 3380 18180 3390 18190
rect 3380 18160 3600 18180
rect 4090 18170 4160 18180
rect 3340 18150 3390 18160
rect 4090 18130 4100 18170
rect 4010 18120 4100 18130
rect 4150 18120 4160 18170
rect 4010 18110 4160 18120
rect 4190 18170 4260 18180
rect 4190 18120 4200 18170
rect 4250 18120 4260 18170
rect 4190 18110 4260 18120
rect 4390 18080 4410 20660
rect 3940 18060 4410 18080
rect 230 15630 640 15640
rect 230 15580 240 15630
rect 290 15620 640 15630
rect 3260 15620 3680 15640
rect 290 15580 300 15620
rect 230 15570 300 15580
rect 3340 15590 3390 15600
rect 3340 15560 3350 15590
rect 3380 15580 3390 15590
rect 3380 15560 3600 15580
rect 4090 15570 4160 15580
rect 3340 15550 3390 15560
rect 4090 15530 4100 15570
rect 4010 15520 4100 15530
rect 4150 15520 4160 15570
rect 4010 15510 4160 15520
rect 4190 15570 4260 15580
rect 4190 15520 4200 15570
rect 4250 15520 4260 15570
rect 4190 15510 4260 15520
rect 4390 15480 4410 18060
rect 7100 16850 7300 21000
rect 6920 16830 7300 16850
rect 3940 15460 4410 15480
rect 4390 13080 4410 15460
rect 6850 14120 6900 14130
rect 6850 14090 6860 14120
rect 6890 14090 6900 14120
rect 6850 14080 6900 14090
rect 6860 13880 6880 14080
rect 6920 13790 6940 14210
rect 6760 13080 6780 13540
rect 6810 13390 6830 13480
rect 6810 13380 6880 13390
rect 6810 13330 6820 13380
rect 6870 13330 6880 13380
rect 6810 13320 6880 13330
rect 6810 13280 6880 13290
rect 6810 13230 6820 13280
rect 6870 13230 6880 13280
rect 6810 13220 6880 13230
rect 4390 13060 6780 13080
rect 230 13030 640 13040
rect 230 12980 240 13030
rect 290 13020 640 13030
rect 3260 13020 3680 13040
rect 290 12980 300 13020
rect 230 12970 300 12980
rect 3340 12990 3390 13000
rect 3340 12960 3350 12990
rect 3380 12980 3390 12990
rect 3380 12960 3600 12980
rect 4090 12970 4160 12980
rect 3340 12950 3390 12960
rect 4090 12930 4100 12970
rect 4010 12920 4100 12930
rect 4150 12920 4160 12970
rect 4010 12910 4160 12920
rect 4190 12970 4260 12980
rect 4190 12920 4200 12970
rect 4250 12920 4260 12970
rect 4190 12910 4260 12920
rect 4390 12880 4410 13060
rect 3940 12860 4410 12880
rect 230 10430 640 10440
rect 230 10380 240 10430
rect 290 10420 640 10430
rect 3260 10420 3680 10440
rect 290 10380 300 10420
rect 230 10370 300 10380
rect 3340 10390 3390 10400
rect 3340 10360 3350 10390
rect 3380 10380 3390 10390
rect 3380 10360 3600 10380
rect 4090 10370 4160 10380
rect 3340 10350 3390 10360
rect 4090 10330 4100 10370
rect 4010 10320 4100 10330
rect 4150 10320 4160 10370
rect 4010 10310 4160 10320
rect 4190 10370 4260 10380
rect 4190 10320 4200 10370
rect 4250 10320 4260 10370
rect 4190 10310 4260 10320
rect 4390 10280 4410 12860
rect 7100 12650 7300 16830
rect 6920 12630 7300 12650
rect 3940 10260 4410 10280
rect 4390 8880 4410 10260
rect 6850 9920 6900 9930
rect 6850 9890 6860 9920
rect 6890 9890 6900 9920
rect 6850 9880 6900 9890
rect 6860 9680 6880 9880
rect 6920 9600 6940 10010
rect 6760 8880 6780 9340
rect 6810 9190 6830 9280
rect 6810 9180 6880 9190
rect 6810 9130 6820 9180
rect 6870 9130 6880 9180
rect 6810 9120 6880 9130
rect 6810 9080 6880 9090
rect 6810 9030 6820 9080
rect 6870 9030 6880 9080
rect 6810 9020 6880 9030
rect 4390 8860 6780 8880
rect 230 7830 640 7840
rect 230 7780 240 7830
rect 290 7820 640 7830
rect 3260 7820 3690 7840
rect 290 7780 300 7820
rect 230 7770 300 7780
rect 3340 7790 3390 7800
rect 3340 7760 3350 7790
rect 3380 7780 3390 7790
rect 3380 7760 3600 7780
rect 4090 7770 4160 7780
rect 3340 7750 3390 7760
rect 4090 7730 4100 7770
rect 4010 7720 4100 7730
rect 4150 7720 4160 7770
rect 4010 7710 4160 7720
rect 4190 7770 4260 7780
rect 4190 7720 4200 7770
rect 4250 7720 4260 7770
rect 4190 7710 4260 7720
rect 4390 7680 4410 8860
rect 7100 8450 7300 12630
rect 6920 8430 7300 8450
rect 3940 7660 4410 7680
rect 230 5230 640 5240
rect 230 5180 240 5230
rect 290 5220 640 5230
rect 3260 5220 3690 5240
rect 290 5180 300 5220
rect 230 5170 300 5180
rect 3340 5190 3390 5200
rect 3340 5160 3350 5190
rect 3380 5180 3390 5190
rect 3380 5160 3610 5180
rect 4090 5170 4160 5180
rect 3340 5150 3390 5160
rect 4090 5130 4100 5170
rect 4010 5120 4100 5130
rect 4150 5120 4160 5170
rect 4010 5110 4160 5120
rect 4190 5170 4260 5180
rect 4190 5120 4200 5170
rect 4250 5120 4260 5170
rect 4190 5110 4260 5120
rect 3940 5080 3980 5090
rect 4390 5080 4410 7660
rect 6850 5720 6900 5730
rect 6850 5690 6860 5720
rect 6890 5690 6900 5720
rect 6850 5680 6900 5690
rect 6860 5480 6880 5680
rect 6920 5390 6940 5810
rect 3940 5060 4410 5080
rect 4390 4680 4410 5060
rect 6760 4680 6780 5140
rect 6810 4990 6830 5080
rect 6810 4980 6880 4990
rect 6810 4930 6820 4980
rect 6870 4930 6880 4980
rect 6810 4920 6880 4930
rect 6810 4880 6880 4890
rect 6810 4830 6820 4880
rect 6870 4830 6880 4880
rect 6810 4820 6880 4830
rect 4390 4660 6780 4680
rect 230 2630 640 2640
rect 230 2580 240 2630
rect 290 2620 640 2630
rect 3260 2620 3690 2640
rect 290 2580 300 2620
rect 3260 2610 3280 2620
rect 3500 2610 3690 2620
rect 230 2570 300 2580
rect 3340 2590 3390 2600
rect 3340 2560 3350 2590
rect 3380 2580 3390 2590
rect 3380 2560 3600 2580
rect 4090 2570 4160 2580
rect 3340 2550 3390 2560
rect 4090 2530 4100 2570
rect 4010 2520 4100 2530
rect 4150 2520 4160 2570
rect 4010 2510 4160 2520
rect 4190 2570 4260 2580
rect 4190 2520 4200 2570
rect 4250 2520 4260 2570
rect 4190 2510 4260 2520
rect 3940 2480 3980 2490
rect 4390 2480 4410 4660
rect 7100 4250 7300 8430
rect 6920 4230 7300 4250
rect 3940 2460 4410 2480
rect 4390 480 4410 2460
rect 6850 1520 6900 1530
rect 6850 1490 6860 1520
rect 6890 1490 6900 1520
rect 6850 1480 6900 1490
rect 6860 1280 6880 1480
rect 6920 1190 6940 1610
rect 6760 480 6780 940
rect 6810 790 6830 880
rect 6810 780 6880 790
rect 6810 730 6820 780
rect 6870 730 6880 780
rect 6810 720 6880 730
rect 6810 680 6880 690
rect 6810 630 6820 680
rect 6870 630 6880 680
rect 6810 620 6880 630
rect 7100 500 7300 4230
rect 7320 13080 7340 16890
rect 9700 16850 9900 21000
rect 9520 16830 9900 16850
rect 9450 14120 9500 14130
rect 9450 14090 9460 14120
rect 9490 14090 9500 14120
rect 9450 14080 9500 14090
rect 9460 13880 9480 14080
rect 9520 13800 9540 14210
rect 9360 13080 9380 13540
rect 9410 13390 9430 13480
rect 9410 13380 9480 13390
rect 9410 13330 9420 13380
rect 9470 13330 9480 13380
rect 9410 13320 9480 13330
rect 9410 13280 9480 13290
rect 9410 13230 9420 13280
rect 9470 13230 9480 13280
rect 9410 13220 9480 13230
rect 7320 13060 9380 13080
rect 7320 8880 7340 13060
rect 9700 12650 9900 16830
rect 9520 12630 9900 12650
rect 9450 9920 9500 9930
rect 9450 9890 9460 9920
rect 9490 9890 9500 9920
rect 9450 9880 9500 9890
rect 9460 9680 9480 9880
rect 9520 9600 9540 10010
rect 9360 8880 9380 9340
rect 9410 9190 9430 9280
rect 9410 9180 9480 9190
rect 9410 9130 9420 9180
rect 9470 9130 9480 9180
rect 9410 9120 9480 9130
rect 9410 9080 9480 9090
rect 9410 9030 9420 9080
rect 9470 9030 9480 9080
rect 9410 9020 9480 9030
rect 7320 8860 9380 8880
rect 7320 4680 7340 8860
rect 9700 8450 9900 12630
rect 9520 8430 9900 8450
rect 9450 5720 9500 5730
rect 9450 5690 9460 5720
rect 9490 5690 9500 5720
rect 9450 5680 9500 5690
rect 9460 5480 9480 5680
rect 9520 5400 9540 5810
rect 9360 4680 9380 5140
rect 9410 4990 9430 5080
rect 9410 4980 9480 4990
rect 9410 4930 9420 4980
rect 9470 4930 9480 4980
rect 9410 4920 9480 4930
rect 9410 4880 9480 4890
rect 9410 4830 9420 4880
rect 9470 4830 9480 4880
rect 9410 4820 9480 4830
rect 7320 4660 9380 4680
rect 4390 460 6780 480
rect 7320 480 7340 4660
rect 9700 4250 9900 8430
rect 9520 4230 9900 4250
rect 9450 1520 9500 1530
rect 9450 1490 9460 1520
rect 9490 1490 9500 1520
rect 9450 1480 9500 1490
rect 9460 1280 9480 1480
rect 9520 1200 9540 1610
rect 9360 480 9380 940
rect 9410 790 9430 880
rect 9410 780 9480 790
rect 9410 730 9420 780
rect 9470 730 9480 780
rect 9410 720 9480 730
rect 9410 680 9480 690
rect 9410 630 9420 680
rect 9470 630 9480 680
rect 9410 620 9480 630
rect 9700 500 9900 4230
rect 7320 460 9380 480
rect 4390 200 4410 460
rect 7320 200 7340 460
rect 4390 190 15250 200
rect 4390 180 15190 190
rect 15180 140 15190 180
rect 15240 140 15250 190
rect 15180 130 15250 140
<< via1 >>
rect 240 20780 290 20830
rect 3350 20760 3380 20790
rect 4100 20720 4150 20770
rect 4200 20720 4250 20770
rect 240 18180 290 18230
rect 3350 18160 3380 18190
rect 4100 18120 4150 18170
rect 4200 18120 4250 18170
rect 240 15580 290 15630
rect 3350 15560 3380 15590
rect 4100 15520 4150 15570
rect 4200 15520 4250 15570
rect 6860 14090 6890 14120
rect 6820 13330 6870 13380
rect 6820 13230 6870 13280
rect 240 12980 290 13030
rect 3350 12960 3380 12990
rect 4100 12920 4150 12970
rect 4200 12920 4250 12970
rect 240 10380 290 10430
rect 3350 10360 3380 10390
rect 4100 10320 4150 10370
rect 4200 10320 4250 10370
rect 6860 9890 6890 9920
rect 6820 9130 6870 9180
rect 6820 9030 6870 9080
rect 240 7780 290 7830
rect 3350 7760 3380 7790
rect 4100 7720 4150 7770
rect 4200 7720 4250 7770
rect 240 5180 290 5230
rect 3350 5160 3380 5190
rect 4100 5120 4150 5170
rect 4200 5120 4250 5170
rect 6860 5690 6890 5720
rect 6820 4930 6870 4980
rect 6820 4830 6870 4880
rect 240 2580 290 2630
rect 3350 2560 3380 2590
rect 4100 2520 4150 2570
rect 4200 2520 4250 2570
rect 6860 1490 6890 1520
rect 6820 730 6870 780
rect 6820 630 6870 680
rect 9460 14090 9490 14120
rect 9420 13330 9470 13380
rect 9420 13230 9470 13280
rect 9460 9890 9490 9920
rect 9420 9130 9470 9180
rect 9420 9030 9470 9080
rect 9460 5690 9490 5720
rect 9420 4930 9470 4980
rect 9420 4830 9470 4880
rect 9460 1490 9490 1520
rect 9420 730 9470 780
rect 9420 630 9470 680
rect 15190 140 15240 190
<< metal2 >>
rect 400 21000 9900 21200
rect 230 20830 300 20840
rect 230 20780 240 20830
rect 290 20780 300 20830
rect 230 20770 300 20780
rect 400 18790 600 21000
rect 4480 20960 4550 20970
rect 4480 20910 4490 20960
rect 4540 20910 4550 20960
rect 4480 20900 4550 20910
rect 4580 20960 4650 20970
rect 4580 20910 4590 20960
rect 4640 20910 4650 20960
rect 4580 20900 4650 20910
rect 4680 20960 4750 20970
rect 4680 20910 4690 20960
rect 4740 20910 4750 20960
rect 4680 20900 4750 20910
rect 4780 20960 4850 20970
rect 4780 20910 4790 20960
rect 4840 20910 4850 20960
rect 4780 20900 4850 20910
rect 4880 20960 4950 20970
rect 4880 20910 4890 20960
rect 4940 20910 4950 20960
rect 4880 20900 4950 20910
rect 4980 20960 5050 20970
rect 4980 20910 4990 20960
rect 5040 20910 5050 20960
rect 4980 20900 5050 20910
rect 5080 20960 5150 20970
rect 5080 20910 5090 20960
rect 5140 20910 5150 20960
rect 5080 20900 5150 20910
rect 5180 20960 5250 20970
rect 5180 20910 5190 20960
rect 5240 20910 5250 20960
rect 5180 20900 5250 20910
rect 3340 20790 3390 20800
rect 3340 20760 3350 20790
rect 3380 20760 3390 20790
rect 3340 20750 3390 20760
rect 4090 20770 4160 20780
rect 4090 20720 4100 20770
rect 4150 20720 4160 20770
rect 4090 20710 4160 20720
rect 4190 20770 4260 20780
rect 4190 20720 4200 20770
rect 4250 20730 4260 20770
rect 4480 20730 4500 20900
rect 4580 20870 4600 20900
rect 4250 20720 4500 20730
rect 4190 20710 4500 20720
rect 4520 20850 4600 20870
rect 400 18740 540 18790
rect 590 18740 630 18790
rect 400 18700 600 18740
rect 230 18230 300 18240
rect 230 18180 240 18230
rect 290 18180 300 18230
rect 230 18170 300 18180
rect 3340 18190 3390 18200
rect 3340 18160 3350 18190
rect 3380 18160 3390 18190
rect 3340 18150 3390 18160
rect 4090 18170 4160 18180
rect 4090 18120 4100 18170
rect 4150 18120 4160 18170
rect 4090 18110 4160 18120
rect 4190 18170 4260 18180
rect 4190 18120 4200 18170
rect 4250 18130 4260 18170
rect 4520 18130 4540 20850
rect 4680 20830 4700 20900
rect 4250 18120 4540 18130
rect 4190 18110 4540 18120
rect 4560 20810 4700 20830
rect 530 16190 600 16200
rect 530 16140 540 16190
rect 590 16140 630 16190
rect 530 16130 600 16140
rect 230 15630 300 15640
rect 230 15580 240 15630
rect 290 15580 300 15630
rect 230 15570 300 15580
rect 3340 15590 3390 15600
rect 3340 15560 3350 15590
rect 3380 15560 3390 15590
rect 3340 15550 3390 15560
rect 4090 15570 4160 15580
rect 4090 15520 4100 15570
rect 4150 15520 4160 15570
rect 4090 15510 4160 15520
rect 4190 15570 4260 15580
rect 4190 15520 4200 15570
rect 4250 15530 4260 15570
rect 4560 15530 4580 20810
rect 4780 20790 4800 20900
rect 4250 15520 4580 15530
rect 4190 15510 4580 15520
rect 4600 20770 4800 20790
rect 530 13590 600 13600
rect 530 13540 540 13590
rect 590 13540 630 13590
rect 530 13530 600 13540
rect 230 13030 300 13040
rect 230 12980 240 13030
rect 290 12980 300 13030
rect 230 12970 300 12980
rect 3340 12990 3390 13000
rect 3340 12960 3350 12990
rect 3380 12960 3390 12990
rect 3340 12950 3390 12960
rect 4090 12970 4160 12980
rect 4090 12920 4100 12970
rect 4150 12920 4160 12970
rect 4090 12910 4160 12920
rect 4190 12970 4260 12980
rect 4190 12920 4200 12970
rect 4250 12930 4260 12970
rect 4600 12930 4620 20770
rect 4880 20750 4900 20900
rect 4250 12920 4620 12930
rect 4190 12910 4620 12920
rect 4640 20730 4900 20750
rect 530 10990 600 11000
rect 530 10940 540 10990
rect 590 10940 630 10990
rect 530 10930 600 10940
rect 230 10430 300 10440
rect 230 10380 240 10430
rect 290 10380 300 10430
rect 230 10370 300 10380
rect 3340 10390 3390 10400
rect 3340 10360 3350 10390
rect 3380 10360 3390 10390
rect 3340 10350 3390 10360
rect 4090 10370 4160 10380
rect 4090 10320 4100 10370
rect 4150 10320 4160 10370
rect 4090 10310 4160 10320
rect 4190 10370 4260 10380
rect 4190 10320 4200 10370
rect 4250 10330 4260 10370
rect 4640 10330 4660 20730
rect 4980 20710 5000 20900
rect 4250 10320 4660 10330
rect 4190 10310 4660 10320
rect 4680 20690 5000 20710
rect 530 8390 600 8400
rect 530 8340 540 8390
rect 590 8340 630 8390
rect 530 8330 600 8340
rect 230 7830 300 7840
rect 230 7780 240 7830
rect 290 7780 300 7830
rect 230 7770 300 7780
rect 3340 7790 3390 7800
rect 3340 7760 3350 7790
rect 3380 7760 3390 7790
rect 3340 7750 3390 7760
rect 4090 7770 4160 7780
rect 4090 7720 4100 7770
rect 4150 7720 4160 7770
rect 4090 7710 4160 7720
rect 4190 7770 4260 7780
rect 4190 7720 4200 7770
rect 4250 7730 4260 7770
rect 4680 7730 4700 20690
rect 5080 20670 5100 20900
rect 4250 7720 4700 7730
rect 4190 7710 4700 7720
rect 4720 20650 5100 20670
rect 530 5790 600 5800
rect 530 5740 540 5790
rect 590 5740 630 5790
rect 530 5730 600 5740
rect 230 5230 300 5240
rect 230 5180 240 5230
rect 290 5180 300 5230
rect 230 5170 300 5180
rect 3340 5190 3390 5200
rect 3340 5160 3350 5190
rect 3380 5160 3390 5190
rect 3340 5150 3390 5160
rect 4090 5170 4160 5180
rect 4090 5120 4100 5170
rect 4150 5120 4160 5170
rect 4090 5110 4160 5120
rect 4190 5170 4260 5180
rect 4190 5120 4200 5170
rect 4250 5130 4260 5170
rect 4720 5130 4740 20650
rect 5180 20630 5200 20900
rect 4250 5120 4740 5130
rect 4190 5110 4740 5120
rect 4760 20610 5200 20630
rect 530 3190 600 3200
rect 530 3140 540 3190
rect 590 3140 630 3190
rect 530 3130 600 3140
rect 230 2630 300 2640
rect 230 2580 240 2630
rect 290 2580 300 2630
rect 230 2570 300 2580
rect 3340 2590 3390 2600
rect 3340 2560 3350 2590
rect 3380 2560 3390 2590
rect 3340 2550 3390 2560
rect 4090 2570 4160 2580
rect 4090 2520 4100 2570
rect 4150 2520 4160 2570
rect 4090 2510 4160 2520
rect 4190 2570 4260 2580
rect 4190 2520 4200 2570
rect 4250 2530 4260 2570
rect 4760 2530 4780 20610
rect 7100 16890 7300 21000
rect 9700 16890 9900 21000
rect 4840 16870 7300 16890
rect 4840 16830 4860 16870
rect 6850 14120 6900 14130
rect 6850 14090 6860 14120
rect 6890 14090 6900 14120
rect 6850 14080 6900 14090
rect 6810 13380 6880 13390
rect 6810 13330 6820 13380
rect 6870 13330 6880 13380
rect 6810 13320 6880 13330
rect 6810 13280 6880 13290
rect 6810 13230 6820 13280
rect 6870 13230 6880 13280
rect 6810 13220 6880 13230
rect 7100 12690 7300 16870
rect 7440 16870 9900 16890
rect 7440 16830 7460 16870
rect 9450 14120 9500 14130
rect 9450 14090 9460 14120
rect 9490 14090 9500 14120
rect 9450 14080 9500 14090
rect 9410 13380 9480 13390
rect 9410 13330 9420 13380
rect 9470 13330 9480 13380
rect 9410 13320 9480 13330
rect 9410 13280 9480 13290
rect 9410 13230 9420 13280
rect 9470 13230 9480 13280
rect 9410 13220 9480 13230
rect 9700 12690 9900 16870
rect 4840 12670 7300 12690
rect 4840 12630 4860 12670
rect 6850 9920 6900 9930
rect 6850 9890 6860 9920
rect 6890 9890 6900 9920
rect 6850 9880 6900 9890
rect 6810 9180 6880 9190
rect 6810 9130 6820 9180
rect 6870 9130 6880 9180
rect 6810 9120 6880 9130
rect 6810 9080 6880 9090
rect 6810 9030 6820 9080
rect 6870 9030 6880 9080
rect 6810 9020 6880 9030
rect 7100 8490 7300 12670
rect 7440 12670 9900 12690
rect 7440 12630 7460 12670
rect 9450 9920 9500 9930
rect 9450 9890 9460 9920
rect 9490 9890 9500 9920
rect 9450 9880 9500 9890
rect 9410 9180 9480 9190
rect 9410 9130 9420 9180
rect 9470 9130 9480 9180
rect 9410 9120 9480 9130
rect 9410 9080 9480 9090
rect 9410 9030 9420 9080
rect 9470 9030 9480 9080
rect 9410 9020 9480 9030
rect 9700 8490 9900 12670
rect 4840 8470 7300 8490
rect 4840 8430 4860 8470
rect 6850 5720 6900 5730
rect 6850 5690 6860 5720
rect 6890 5690 6900 5720
rect 6850 5680 6900 5690
rect 6810 4980 6880 4990
rect 6810 4930 6820 4980
rect 6870 4930 6880 4980
rect 6810 4920 6880 4930
rect 6810 4880 6880 4890
rect 6810 4830 6820 4880
rect 6870 4830 6880 4880
rect 6810 4820 6880 4830
rect 7100 4290 7300 8470
rect 7440 8470 9900 8490
rect 7440 8430 7460 8470
rect 9450 5720 9500 5730
rect 9450 5690 9460 5720
rect 9490 5690 9500 5720
rect 9450 5680 9500 5690
rect 9410 4980 9480 4990
rect 9410 4930 9420 4980
rect 9470 4930 9480 4980
rect 9410 4920 9480 4930
rect 9410 4880 9480 4890
rect 9410 4830 9420 4880
rect 9470 4830 9480 4880
rect 9410 4820 9480 4830
rect 9700 4290 9900 8470
rect 4840 4270 7300 4290
rect 4840 4230 4860 4270
rect 4250 2520 4780 2530
rect 4190 2510 4780 2520
rect 6850 1520 6900 1530
rect 6850 1490 6860 1520
rect 6890 1490 6900 1520
rect 6850 1480 6900 1490
rect 6810 780 6880 790
rect 6810 730 6820 780
rect 6870 730 6880 780
rect 6810 720 6880 730
rect 6810 680 6880 690
rect 6810 630 6820 680
rect 6870 630 6880 680
rect 6810 620 6880 630
rect 530 590 600 600
rect 530 540 540 590
rect 590 540 630 590
rect 530 530 600 540
rect 7100 500 7300 4270
rect 7440 4270 9900 4290
rect 7440 4230 7460 4270
rect 9450 1520 9500 1530
rect 9450 1490 9460 1520
rect 9490 1490 9500 1520
rect 9450 1480 9500 1490
rect 9410 780 9480 790
rect 9410 730 9420 780
rect 9470 730 9480 780
rect 9410 720 9480 730
rect 9410 680 9480 690
rect 9410 630 9420 680
rect 9470 630 9480 680
rect 9410 620 9480 630
rect 9700 500 9900 4270
rect 15180 190 15250 200
rect 15180 140 15190 190
rect 15240 140 15250 190
rect 15180 130 15250 140
<< via2 >>
rect 240 20780 290 20830
rect 4490 20910 4540 20960
rect 4590 20910 4640 20960
rect 4690 20910 4740 20960
rect 4790 20910 4840 20960
rect 4890 20910 4940 20960
rect 4990 20910 5040 20960
rect 5090 20910 5140 20960
rect 5190 20910 5240 20960
rect 4100 20720 4150 20770
rect 4200 20720 4250 20770
rect 540 18740 590 18790
rect 240 18180 290 18230
rect 4100 18120 4150 18170
rect 4200 18120 4250 18170
rect 540 16140 590 16190
rect 240 15580 290 15630
rect 4100 15520 4150 15570
rect 4200 15520 4250 15570
rect 540 13540 590 13590
rect 240 12980 290 13030
rect 4100 12920 4150 12970
rect 4200 12920 4250 12970
rect 540 10940 590 10990
rect 240 10380 290 10430
rect 4100 10320 4150 10370
rect 4200 10320 4250 10370
rect 540 8340 590 8390
rect 240 7780 290 7830
rect 4100 7720 4150 7770
rect 4200 7720 4250 7770
rect 540 5740 590 5790
rect 240 5180 290 5230
rect 4100 5120 4150 5170
rect 4200 5120 4250 5170
rect 540 3140 590 3190
rect 240 2580 290 2630
rect 4100 2520 4150 2570
rect 4200 2520 4250 2570
rect 6820 13330 6870 13380
rect 6820 13230 6870 13280
rect 9420 13330 9470 13380
rect 9420 13230 9470 13280
rect 6820 9130 6870 9180
rect 6820 9030 6870 9080
rect 9420 9130 9470 9180
rect 9420 9030 9470 9080
rect 6820 4930 6870 4980
rect 6820 4830 6870 4880
rect 9420 4930 9470 4980
rect 9420 4830 9470 4880
rect 6820 730 6870 780
rect 6820 630 6870 680
rect 540 540 590 590
rect 9420 730 9470 780
rect 9420 630 9470 680
rect 15190 140 15240 190
<< metal3 >>
rect 9680 22430 9750 22440
rect 9680 22380 9690 22430
rect 9740 22380 9750 22430
rect 9680 22370 9750 22380
rect 9960 22430 10030 22440
rect 9960 22380 9970 22430
rect 10020 22380 10030 22430
rect 9960 22370 10030 22380
rect 10230 22430 10300 22440
rect 10230 22380 10240 22430
rect 10290 22380 10300 22430
rect 10230 22370 10300 22380
rect 10510 22430 10580 22440
rect 10510 22380 10520 22430
rect 10570 22380 10580 22430
rect 10510 22370 10580 22380
rect 10790 22430 10860 22440
rect 10790 22380 10800 22430
rect 10850 22380 10860 22430
rect 10790 22370 10860 22380
rect 11070 22430 11140 22440
rect 11070 22380 11080 22430
rect 11130 22380 11140 22430
rect 11070 22370 11140 22380
rect 11340 22430 11410 22440
rect 11340 22380 11350 22430
rect 11400 22380 11410 22430
rect 11340 22370 11410 22380
rect 11610 22430 11680 22440
rect 11610 22380 11620 22430
rect 11670 22380 11680 22430
rect 11610 22370 11680 22380
rect 11890 22430 11960 22440
rect 11890 22380 11900 22430
rect 11950 22380 11960 22430
rect 11890 22370 11960 22380
rect 12170 22430 12240 22440
rect 12170 22380 12180 22430
rect 12230 22380 12240 22430
rect 12170 22370 12240 22380
rect 12450 22430 12520 22440
rect 12450 22380 12460 22430
rect 12510 22380 12520 22430
rect 12450 22370 12520 22380
rect 12720 22430 12790 22440
rect 12720 22380 12730 22430
rect 12780 22380 12790 22430
rect 12720 22370 12790 22380
rect 13000 22430 13070 22440
rect 13000 22380 13010 22430
rect 13060 22380 13070 22430
rect 13000 22370 13070 22380
rect 13280 22430 13350 22440
rect 13280 22380 13290 22430
rect 13340 22380 13350 22430
rect 13280 22370 13350 22380
rect 13550 22430 13620 22440
rect 13550 22380 13560 22430
rect 13610 22380 13620 22430
rect 13550 22370 13620 22380
rect 13830 22430 13900 22440
rect 13830 22380 13840 22430
rect 13890 22380 13900 22430
rect 13830 22370 13900 22380
rect 9680 22100 9710 22370
rect 9960 22100 9990 22370
rect 10230 22100 10260 22370
rect 10510 22100 10540 22370
rect 9680 22090 9750 22100
rect 9680 22040 9690 22090
rect 9740 22040 9750 22090
rect 9680 22030 9750 22040
rect 9960 22090 10030 22100
rect 9960 22040 9970 22090
rect 10020 22040 10030 22090
rect 9960 22030 10030 22040
rect 10230 22090 10300 22100
rect 10230 22040 10240 22090
rect 10290 22040 10300 22090
rect 10230 22030 10300 22040
rect 10510 22090 10580 22100
rect 10510 22040 10520 22090
rect 10570 22040 10580 22090
rect 10510 22030 10580 22040
rect 11900 21670 11930 22370
rect 4480 21640 11930 21670
rect 4480 20960 4510 21640
rect 12180 21610 12210 22370
rect 4580 21580 12210 21610
rect 4480 20940 4490 20960
rect 4580 20960 4610 21580
rect 12450 21550 12480 22370
rect 4680 21520 12480 21550
rect 4580 20940 4590 20960
rect 4680 20960 4710 21520
rect 12730 21490 12760 22370
rect 4780 21460 12760 21490
rect 4680 20940 4690 20960
rect 4780 20960 4810 21460
rect 13010 21430 13040 22370
rect 4880 21400 13040 21430
rect 4780 20940 4790 20960
rect 4880 20960 4910 21400
rect 13290 21370 13320 22370
rect 4980 21340 13320 21370
rect 4880 20940 4890 20960
rect 4980 20960 5010 21340
rect 13560 21310 13590 22370
rect 5080 21280 13590 21310
rect 4980 20940 4990 20960
rect 5080 20960 5130 21280
rect 13830 21250 13860 22370
rect 5180 21220 13860 21250
rect 5080 20940 5090 20960
rect 5180 20960 5210 21220
rect 5180 20940 5190 20960
rect 230 20830 300 20840
rect 230 20780 240 20830
rect 290 20780 300 20830
rect 230 20770 300 20780
rect 4090 20770 4160 20780
rect 4090 20720 4100 20770
rect 4150 20720 4160 20770
rect 4090 20710 4160 20720
rect 4190 20770 4260 20780
rect 4190 20720 4200 20770
rect 4250 20720 4260 20770
rect 4190 20710 4260 20720
rect 530 18790 600 18800
rect 530 18740 540 18790
rect 590 18740 600 18790
rect 530 18730 600 18740
rect 230 18230 300 18240
rect 230 18180 240 18230
rect 290 18180 300 18230
rect 230 18170 300 18180
rect 4090 18170 4160 18180
rect 4090 18120 4100 18170
rect 4150 18120 4160 18170
rect 4090 18110 4160 18120
rect 4190 18170 4260 18180
rect 4190 18120 4200 18170
rect 4250 18120 4260 18170
rect 4190 18110 4260 18120
rect 530 16190 600 16200
rect 530 16140 540 16190
rect 590 16140 600 16190
rect 530 16130 600 16140
rect 230 15630 300 15640
rect 230 15580 240 15630
rect 290 15580 300 15630
rect 230 15570 300 15580
rect 4090 15570 4160 15580
rect 4090 15520 4100 15570
rect 4150 15520 4160 15570
rect 4090 15510 4160 15520
rect 4190 15570 4260 15580
rect 4190 15520 4200 15570
rect 4250 15520 4260 15570
rect 4190 15510 4260 15520
rect 530 13590 600 13600
rect 530 13540 540 13590
rect 590 13540 600 13590
rect 530 13530 600 13540
rect 6810 13380 6880 13390
rect 6810 13330 6820 13380
rect 6870 13330 6880 13380
rect 6810 13320 6880 13330
rect 9410 13380 9480 13390
rect 9410 13330 9420 13380
rect 9470 13330 9480 13380
rect 9410 13320 9480 13330
rect 6810 13280 6880 13290
rect 6810 13230 6820 13280
rect 6870 13230 6880 13280
rect 6810 13220 6880 13230
rect 9410 13280 9480 13290
rect 9410 13230 9420 13280
rect 9470 13230 9480 13280
rect 9410 13220 9480 13230
rect 230 13030 300 13040
rect 230 12980 240 13030
rect 290 12980 300 13030
rect 230 12970 300 12980
rect 4090 12970 4160 12980
rect 4090 12920 4100 12970
rect 4150 12920 4160 12970
rect 4090 12910 4160 12920
rect 4190 12970 4260 12980
rect 4190 12920 4200 12970
rect 4250 12920 4260 12970
rect 4190 12910 4260 12920
rect 530 10990 600 11000
rect 530 10940 540 10990
rect 590 10940 600 10990
rect 530 10930 600 10940
rect 230 10430 300 10440
rect 230 10380 240 10430
rect 290 10380 300 10430
rect 230 10370 300 10380
rect 4090 10370 4160 10380
rect 4090 10320 4100 10370
rect 4150 10320 4160 10370
rect 4090 10310 4160 10320
rect 4190 10370 4260 10380
rect 4190 10320 4200 10370
rect 4250 10320 4260 10370
rect 4190 10310 4260 10320
rect 6810 9180 6880 9190
rect 6810 9130 6820 9180
rect 6870 9130 6880 9180
rect 6810 9120 6880 9130
rect 9410 9180 9480 9190
rect 9410 9130 9420 9180
rect 9470 9130 9480 9180
rect 9410 9120 9480 9130
rect 6810 9080 6880 9090
rect 6810 9030 6820 9080
rect 6870 9030 6880 9080
rect 6810 9020 6880 9030
rect 9410 9080 9480 9090
rect 9410 9030 9420 9080
rect 9470 9030 9480 9080
rect 9410 9020 9480 9030
rect 530 8390 600 8400
rect 530 8340 540 8390
rect 590 8340 600 8390
rect 530 8330 600 8340
rect 230 7830 300 7840
rect 230 7780 240 7830
rect 290 7780 300 7830
rect 230 7770 300 7780
rect 4090 7770 4160 7780
rect 4090 7720 4100 7770
rect 4150 7720 4160 7770
rect 4090 7710 4160 7720
rect 4190 7770 4260 7780
rect 4190 7720 4200 7770
rect 4250 7720 4260 7770
rect 4190 7710 4260 7720
rect 530 5790 600 5800
rect 530 5740 540 5790
rect 590 5740 600 5790
rect 530 5730 600 5740
rect 230 5230 300 5240
rect 230 5180 240 5230
rect 290 5180 300 5230
rect 230 5170 300 5180
rect 4090 5170 4160 5180
rect 4090 5120 4100 5170
rect 4150 5120 4160 5170
rect 4090 5110 4160 5120
rect 4190 5170 4260 5180
rect 4190 5120 4200 5170
rect 4250 5120 4260 5170
rect 4190 5110 4260 5120
rect 6810 4980 6880 4990
rect 6810 4930 6820 4980
rect 6870 4930 6880 4980
rect 6810 4920 6880 4930
rect 9410 4980 9480 4990
rect 9410 4930 9420 4980
rect 9470 4930 9480 4980
rect 9410 4920 9480 4930
rect 6810 4880 6880 4890
rect 6810 4830 6820 4880
rect 6870 4830 6880 4880
rect 6810 4820 6880 4830
rect 9410 4880 9480 4890
rect 9410 4830 9420 4880
rect 9470 4830 9480 4880
rect 9410 4820 9480 4830
rect 530 3190 600 3200
rect 530 3140 540 3190
rect 590 3140 600 3190
rect 530 3130 600 3140
rect 230 2630 300 2640
rect 230 2580 240 2630
rect 290 2580 300 2630
rect 230 2570 300 2580
rect 4090 2570 4160 2580
rect 4090 2520 4100 2570
rect 4150 2520 4160 2570
rect 4090 2510 4160 2520
rect 4190 2570 4260 2580
rect 4190 2520 4200 2570
rect 4250 2520 4260 2570
rect 4190 2510 4260 2520
rect 6810 780 6880 790
rect 6810 730 6820 780
rect 6870 730 6880 780
rect 6810 720 6880 730
rect 9410 780 9480 790
rect 9410 730 9420 780
rect 9470 730 9480 780
rect 9410 720 9480 730
rect 6810 680 6880 690
rect 6810 630 6820 680
rect 6870 630 6880 680
rect 6810 620 6880 630
rect 9410 680 9480 690
rect 9410 630 9420 680
rect 9470 630 9480 680
rect 9410 620 9480 630
rect 530 590 600 600
rect 530 540 540 590
rect 590 540 600 590
rect 530 530 600 540
rect 15180 190 15250 200
rect 15180 140 15190 190
rect 15240 140 15250 190
rect 15180 130 15250 140
<< rmetal3 >>
rect 4510 20960 4550 20970
rect 4480 20910 4490 20940
rect 4540 20910 4550 20960
rect 4480 20900 4550 20910
rect 4610 20960 4650 20970
rect 4580 20910 4590 20940
rect 4640 20910 4650 20960
rect 4580 20900 4650 20910
rect 4710 20960 4750 20970
rect 4680 20910 4690 20940
rect 4740 20910 4750 20960
rect 4680 20900 4750 20910
rect 4810 20960 4850 20970
rect 4780 20910 4790 20940
rect 4840 20910 4850 20960
rect 4780 20900 4850 20910
rect 4910 20960 4950 20970
rect 4880 20910 4890 20940
rect 4940 20910 4950 20960
rect 4880 20900 4950 20910
rect 5010 20960 5050 20970
rect 4980 20910 4990 20940
rect 5040 20910 5050 20960
rect 4980 20900 5050 20910
rect 5130 20960 5150 20970
rect 5080 20910 5090 20940
rect 5140 20910 5150 20960
rect 5080 20900 5150 20910
rect 5210 20960 5250 20970
rect 5180 20910 5190 20940
rect 5240 20910 5250 20960
rect 5180 20900 5250 20910
<< via3 >>
rect 9690 22380 9740 22430
rect 9970 22380 10020 22430
rect 10240 22380 10290 22430
rect 10520 22380 10570 22430
rect 10800 22380 10850 22430
rect 11080 22380 11130 22430
rect 11350 22380 11400 22430
rect 11620 22380 11670 22430
rect 11900 22380 11950 22430
rect 12180 22380 12230 22430
rect 12460 22380 12510 22430
rect 12730 22380 12780 22430
rect 13010 22380 13060 22430
rect 13290 22380 13340 22430
rect 13560 22380 13610 22430
rect 13840 22380 13890 22430
rect 9690 22040 9740 22090
rect 9970 22040 10020 22090
rect 10240 22040 10290 22090
rect 10520 22040 10570 22090
rect 240 20780 290 20830
rect 4100 20720 4150 20770
rect 4200 20720 4250 20770
rect 540 18740 590 18790
rect 240 18180 290 18230
rect 4100 18120 4150 18170
rect 4200 18120 4250 18170
rect 540 16140 590 16190
rect 240 15580 290 15630
rect 4100 15520 4150 15570
rect 4200 15520 4250 15570
rect 540 13540 590 13590
rect 6820 13330 6870 13380
rect 9420 13330 9470 13380
rect 6820 13230 6870 13280
rect 9420 13230 9470 13280
rect 240 12980 290 13030
rect 4100 12920 4150 12970
rect 4200 12920 4250 12970
rect 540 10940 590 10990
rect 240 10380 290 10430
rect 4100 10320 4150 10370
rect 4200 10320 4250 10370
rect 6820 9130 6870 9180
rect 9420 9130 9470 9180
rect 6820 9030 6870 9080
rect 9420 9030 9470 9080
rect 540 8340 590 8390
rect 240 7780 290 7830
rect 4100 7720 4150 7770
rect 4200 7720 4250 7770
rect 540 5740 590 5790
rect 240 5180 290 5230
rect 4100 5120 4150 5170
rect 4200 5120 4250 5170
rect 6820 4930 6870 4980
rect 9420 4930 9470 4980
rect 6820 4830 6870 4880
rect 9420 4830 9470 4880
rect 540 3140 590 3190
rect 240 2580 290 2630
rect 4100 2520 4150 2570
rect 4200 2520 4250 2570
rect 6820 730 6870 780
rect 9420 730 9470 780
rect 6820 630 6870 680
rect 9420 630 9470 680
rect 540 540 590 590
rect 15190 140 15240 190
<< metal4 >>
rect 3067 22510 3097 22576
rect 3343 22510 3373 22576
rect 3619 22510 3649 22576
rect 3895 22510 3925 22576
rect 4171 22510 4201 22576
rect 3067 22476 3100 22510
rect 3343 22476 3380 22510
rect 3619 22476 3650 22510
rect 3895 22476 3930 22510
rect 3070 22440 3100 22476
rect 3350 22440 3380 22476
rect 3620 22440 3650 22476
rect 3900 22440 3930 22476
rect 4170 22476 4201 22510
rect 4447 22510 4477 22576
rect 4723 22510 4753 22576
rect 4999 22510 5029 22576
rect 5275 22510 5305 22576
rect 5551 22510 5581 22576
rect 4447 22476 4480 22510
rect 4723 22476 4760 22510
rect 4999 22476 5030 22510
rect 5275 22476 5310 22510
rect 4170 22440 4200 22476
rect 4450 22440 4480 22476
rect 4730 22440 4760 22476
rect 5000 22440 5030 22476
rect 5280 22440 5310 22476
rect 5550 22476 5581 22510
rect 5827 22510 5857 22576
rect 6103 22510 6133 22576
rect 6379 22510 6409 22576
rect 6655 22510 6685 22576
rect 6931 22510 6961 22576
rect 5827 22476 5860 22510
rect 6103 22476 6140 22510
rect 6379 22476 6410 22510
rect 6655 22476 6690 22510
rect 5550 22440 5580 22476
rect 5830 22440 5860 22476
rect 6110 22440 6140 22476
rect 6380 22440 6410 22476
rect 6660 22440 6690 22476
rect 6930 22476 6961 22510
rect 7207 22510 7237 22576
rect 7483 22510 7513 22576
rect 7759 22510 7789 22576
rect 8035 22510 8065 22576
rect 8311 22510 8341 22576
rect 7207 22476 7240 22510
rect 7483 22476 7520 22510
rect 7759 22476 7790 22510
rect 8035 22476 8070 22510
rect 6930 22440 6960 22476
rect 7210 22440 7240 22476
rect 7490 22440 7520 22476
rect 7760 22440 7790 22476
rect 8040 22440 8070 22476
rect 8310 22476 8341 22510
rect 8587 22510 8617 22576
rect 8863 22510 8893 22576
rect 8587 22476 8620 22510
rect 8310 22440 8340 22476
rect 8590 22440 8620 22476
rect 8860 22476 8893 22510
rect 9139 22510 9169 22576
rect 9415 22510 9445 22576
rect 9139 22476 9170 22510
rect 9415 22476 9450 22510
rect 9691 22490 9721 22576
rect 8860 22440 8890 22476
rect 9140 22440 9170 22476
rect 9420 22440 9450 22476
rect 9690 22476 9721 22490
rect 9967 22490 9997 22576
rect 10243 22490 10273 22576
rect 9967 22476 10000 22490
rect 9690 22440 9720 22476
rect 9970 22440 10000 22476
rect 10240 22476 10273 22490
rect 10519 22490 10549 22576
rect 10795 22490 10825 22576
rect 11071 22490 11101 22576
rect 10519 22476 10550 22490
rect 10240 22440 10270 22476
rect 10520 22440 10550 22476
rect 10790 22440 10830 22490
rect 11070 22476 11101 22490
rect 11347 22500 11377 22576
rect 11623 22500 11653 22576
rect 11899 22500 11929 22576
rect 12175 22500 12205 22576
rect 12451 22500 12481 22576
rect 12727 22500 12757 22576
rect 13003 22500 13033 22576
rect 11347 22476 11380 22500
rect 11070 22440 11100 22476
rect 11350 22440 11380 22476
rect 11620 22476 11653 22500
rect 11890 22476 11929 22500
rect 12170 22476 12205 22500
rect 12450 22476 12481 22500
rect 12720 22476 12757 22500
rect 13000 22476 13033 22500
rect 13279 22500 13309 22576
rect 13555 22500 13585 22576
rect 13831 22500 13861 22576
rect 13279 22476 13310 22500
rect 11620 22440 11650 22476
rect 11890 22440 11920 22476
rect 12170 22440 12200 22476
rect 12450 22440 12480 22476
rect 12720 22440 12750 22476
rect 13000 22440 13030 22476
rect 13280 22440 13310 22476
rect 13550 22476 13585 22500
rect 13830 22476 13861 22500
rect 14107 22476 14137 22576
rect 14383 22476 14413 22576
rect 14659 22476 14689 22576
rect 13550 22440 13580 22476
rect 13830 22440 13860 22476
rect 630 22410 9450 22440
rect 9680 22430 9750 22440
rect 630 22080 660 22410
rect 9680 22380 9690 22430
rect 9740 22380 9750 22430
rect 9680 22370 9750 22380
rect 9960 22430 10030 22440
rect 9960 22380 9970 22430
rect 10020 22380 10030 22430
rect 9960 22370 10030 22380
rect 10230 22430 10300 22440
rect 10230 22380 10240 22430
rect 10290 22380 10300 22430
rect 10230 22370 10300 22380
rect 10510 22430 10580 22440
rect 10510 22380 10520 22430
rect 10570 22380 10580 22430
rect 10510 22370 10580 22380
rect 10790 22430 10860 22440
rect 10790 22380 10800 22430
rect 10850 22380 10860 22430
rect 10790 22370 10860 22380
rect 11070 22430 11140 22440
rect 11070 22380 11080 22430
rect 11130 22380 11140 22430
rect 11070 22370 11140 22380
rect 11340 22430 11410 22440
rect 11340 22380 11350 22430
rect 11400 22380 11410 22430
rect 11340 22370 11410 22380
rect 11610 22430 11680 22440
rect 11610 22380 11620 22430
rect 11670 22380 11680 22430
rect 11610 22370 11680 22380
rect 11890 22430 11960 22440
rect 11890 22380 11900 22430
rect 11950 22380 11960 22430
rect 11890 22370 11960 22380
rect 12170 22430 12240 22440
rect 12170 22380 12180 22430
rect 12230 22380 12240 22430
rect 12170 22370 12240 22380
rect 12450 22430 12520 22440
rect 12450 22380 12460 22430
rect 12510 22380 12520 22430
rect 12450 22370 12520 22380
rect 12720 22430 12790 22440
rect 12720 22380 12730 22430
rect 12780 22380 12790 22430
rect 12720 22370 12790 22380
rect 13000 22430 13070 22440
rect 13000 22380 13010 22430
rect 13060 22380 13070 22430
rect 13000 22370 13070 22380
rect 13280 22430 13350 22440
rect 13280 22380 13290 22430
rect 13340 22380 13350 22430
rect 13280 22370 13350 22380
rect 13550 22430 13620 22440
rect 13550 22380 13560 22430
rect 13610 22380 13620 22430
rect 13550 22370 13620 22380
rect 13830 22430 13900 22440
rect 13830 22380 13840 22430
rect 13890 22380 13900 22430
rect 13830 22370 13900 22380
rect 10790 22340 10820 22370
rect 570 22076 660 22080
rect 100 20830 300 22076
rect 100 20780 240 20830
rect 290 20780 300 20830
rect 100 18230 300 20780
rect 100 18180 240 18230
rect 290 18180 300 18230
rect 100 15630 300 18180
rect 100 15580 240 15630
rect 290 15580 300 15630
rect 100 13030 300 15580
rect 100 12980 240 13030
rect 290 12980 300 13030
rect 100 10430 300 12980
rect 100 10380 240 10430
rect 290 10380 300 10430
rect 100 7830 300 10380
rect 100 7780 240 7830
rect 290 7780 300 7830
rect 100 5230 300 7780
rect 100 5180 240 5230
rect 290 5180 300 5230
rect 100 2630 300 5180
rect 100 2580 240 2630
rect 290 2580 300 2630
rect 100 500 300 2580
rect 400 22050 660 22076
rect 7090 22310 10820 22340
rect 400 18790 600 22050
rect 4090 20770 4160 20780
rect 4090 20720 4100 20770
rect 4150 20740 4160 20770
rect 4190 20770 4260 20780
rect 4190 20740 4200 20770
rect 4150 20720 4200 20740
rect 4250 20720 4260 20770
rect 4090 20710 4260 20720
rect 400 18740 540 18790
rect 590 18740 600 18790
rect 400 16190 600 18740
rect 4090 18170 4160 18180
rect 4090 18120 4100 18170
rect 4150 18140 4160 18170
rect 4190 18170 4260 18180
rect 4190 18140 4200 18170
rect 4150 18120 4200 18140
rect 4250 18120 4260 18170
rect 4090 18110 4260 18120
rect 400 16140 540 16190
rect 590 16140 600 16190
rect 400 13590 600 16140
rect 4090 15570 4160 15580
rect 4090 15520 4100 15570
rect 4150 15540 4160 15570
rect 4190 15570 4260 15580
rect 4190 15540 4200 15570
rect 4150 15520 4200 15540
rect 4250 15520 4260 15570
rect 4090 15510 4260 15520
rect 400 13540 540 13590
rect 590 13540 600 13590
rect 400 10990 600 13540
rect 6810 13380 6880 13390
rect 6810 13330 6820 13380
rect 6870 13330 6880 13380
rect 6810 13320 6880 13330
rect 6810 13290 6840 13320
rect 6810 13280 6880 13290
rect 6810 13230 6820 13280
rect 6870 13250 6880 13280
rect 7090 13250 7120 22310
rect 11070 22280 11100 22370
rect 6870 13230 7120 13250
rect 6810 13220 7120 13230
rect 7150 22250 11100 22280
rect 4090 12970 4160 12980
rect 4090 12920 4100 12970
rect 4150 12940 4160 12970
rect 4190 12970 4260 12980
rect 4190 12940 4200 12970
rect 4150 12920 4200 12940
rect 4250 12920 4260 12970
rect 4090 12910 4260 12920
rect 400 10940 540 10990
rect 590 10940 600 10990
rect 400 8390 600 10940
rect 4090 10370 4160 10380
rect 4090 10320 4100 10370
rect 4150 10340 4160 10370
rect 4190 10370 4260 10380
rect 4190 10340 4200 10370
rect 4150 10320 4200 10340
rect 4250 10320 4260 10370
rect 4090 10310 4260 10320
rect 6810 9180 6880 9190
rect 6810 9130 6820 9180
rect 6870 9130 6880 9180
rect 6810 9120 6880 9130
rect 6810 9090 6840 9120
rect 6810 9080 6880 9090
rect 6810 9030 6820 9080
rect 6870 9050 6880 9080
rect 7150 9050 7180 22250
rect 11340 22220 11370 22370
rect 6870 9030 7180 9050
rect 6810 9020 7180 9030
rect 7210 22190 11370 22220
rect 400 8340 540 8390
rect 590 8340 600 8390
rect 400 5790 600 8340
rect 4090 7770 4160 7780
rect 4090 7720 4100 7770
rect 4150 7740 4160 7770
rect 4190 7770 4260 7780
rect 4190 7740 4200 7770
rect 4150 7720 4200 7740
rect 4250 7720 4260 7770
rect 4090 7710 4260 7720
rect 400 5740 540 5790
rect 590 5740 600 5790
rect 400 3190 600 5740
rect 4090 5170 4160 5180
rect 4090 5120 4100 5170
rect 4150 5140 4160 5170
rect 4190 5170 4260 5180
rect 4190 5140 4200 5170
rect 4150 5120 4200 5140
rect 4250 5120 4260 5170
rect 4090 5110 4260 5120
rect 6810 4980 6880 4990
rect 6810 4930 6820 4980
rect 6870 4930 6880 4980
rect 6810 4920 6880 4930
rect 6810 4890 6840 4920
rect 6810 4880 6880 4890
rect 6810 4830 6820 4880
rect 6870 4850 6880 4880
rect 7210 4850 7240 22190
rect 11610 22160 11640 22370
rect 6870 4830 7240 4850
rect 6810 4820 7240 4830
rect 7270 22130 11640 22160
rect 400 3140 540 3190
rect 590 3140 600 3190
rect 400 590 600 3140
rect 4090 2570 4160 2580
rect 4090 2520 4100 2570
rect 4150 2540 4160 2570
rect 4190 2570 4260 2580
rect 4190 2540 4200 2570
rect 4150 2520 4200 2540
rect 4250 2520 4260 2570
rect 4090 2510 4260 2520
rect 6810 780 6880 790
rect 6810 730 6820 780
rect 6870 730 6880 780
rect 6810 720 6880 730
rect 6810 690 6840 720
rect 6810 680 6880 690
rect 6810 630 6820 680
rect 6870 650 6880 680
rect 7270 650 7300 22130
rect 9680 22090 9750 22100
rect 9680 22040 9690 22090
rect 9740 22040 9750 22090
rect 9680 22030 9750 22040
rect 9960 22090 10030 22100
rect 9960 22040 9970 22090
rect 10020 22040 10030 22090
rect 9960 22030 10030 22040
rect 10230 22090 10300 22100
rect 10230 22040 10240 22090
rect 10290 22040 10300 22090
rect 10230 22030 10300 22040
rect 10510 22090 10580 22100
rect 10510 22040 10520 22090
rect 10570 22040 10580 22090
rect 10510 22030 10580 22040
rect 9410 13380 9480 13390
rect 9410 13330 9420 13380
rect 9470 13330 9480 13380
rect 9410 13320 9480 13330
rect 9410 13290 9440 13320
rect 9410 13280 9480 13290
rect 9410 13230 9420 13280
rect 9470 13250 9480 13280
rect 9690 13250 9720 22030
rect 9960 22000 9990 22030
rect 9470 13230 9720 13250
rect 9410 13220 9720 13230
rect 9750 21970 9990 22000
rect 9410 9180 9480 9190
rect 9410 9130 9420 9180
rect 9470 9130 9480 9180
rect 9410 9120 9480 9130
rect 9410 9090 9440 9120
rect 9410 9080 9480 9090
rect 9410 9030 9420 9080
rect 9470 9050 9480 9080
rect 9750 9050 9780 21970
rect 10230 21940 10260 22030
rect 9470 9030 9780 9050
rect 9410 9020 9780 9030
rect 9810 21910 10260 21940
rect 9410 4980 9480 4990
rect 9410 4930 9420 4980
rect 9470 4930 9480 4980
rect 9410 4920 9480 4930
rect 9410 4890 9440 4920
rect 9410 4880 9480 4890
rect 9410 4830 9420 4880
rect 9470 4850 9480 4880
rect 9810 4850 9840 21910
rect 10510 21880 10540 22030
rect 9470 4830 9840 4850
rect 9410 4820 9840 4830
rect 9870 21850 10540 21880
rect 6870 630 7300 650
rect 6810 620 7300 630
rect 9410 780 9480 790
rect 9410 730 9420 780
rect 9470 730 9480 780
rect 9410 720 9480 730
rect 9410 690 9440 720
rect 9410 680 9480 690
rect 9410 630 9420 680
rect 9470 650 9480 680
rect 9870 650 9900 21850
rect 9470 630 9900 650
rect 9410 620 9900 630
rect 400 540 540 590
rect 590 540 600 590
rect 400 500 600 540
rect 15180 190 15250 200
rect 15180 140 15190 190
rect 15240 140 15250 190
rect 15180 130 15250 140
rect 15180 100 15210 130
rect 1657 0 1747 100
rect 3589 0 3679 100
rect 5521 0 5611 100
rect 7453 0 7543 100
rect 9385 0 9475 100
rect 11317 0 11407 100
rect 13249 0 13339 100
rect 15180 70 15271 100
rect 15181 0 15271 70
use bias_generator  bias_generator_0 bias_generator/mag
timestamp 1722981971
transform 1 0 -978 0 1 -680
box 1578 1180 5350 3320
use bias_generator  bias_generator_1
timestamp 1722981971
transform 1 0 -978 0 1 1920
box 1578 1180 5350 3320
use bias_generator  bias_generator_2
timestamp 1722981971
transform 1 0 -978 0 1 4520
box 1578 1180 5350 3320
use bias_generator  bias_generator_3
timestamp 1722981971
transform 1 0 -978 0 1 7120
box 1578 1180 5350 3320
use bias_generator  bias_generator_4
timestamp 1722981971
transform 1 0 -978 0 1 9720
box 1578 1180 5350 3320
use bias_generator  bias_generator_5
timestamp 1722981971
transform 1 0 -978 0 1 12320
box 1578 1180 5350 3320
use bias_generator  bias_generator_6
timestamp 1722981971
transform 1 0 -978 0 1 14920
box 1578 1180 5350 3320
use bias_generator  bias_generator_7
timestamp 1722981971
transform 1 0 -978 0 1 17520
box 1578 1180 5350 3320
use bias_generator  bias_generator_8
timestamp 1722981971
transform 0 1 3620 -1 0 5850
box 1578 1180 5350 3320
use bias_generator  bias_generator_9
timestamp 1722981971
transform 0 1 3620 -1 0 10050
box 1578 1180 5350 3320
use bias_generator  bias_generator_10
timestamp 1722981971
transform 0 1 3620 -1 0 14250
box 1578 1180 5350 3320
use bias_generator  bias_generator_11
timestamp 1722981971
transform 0 1 3620 -1 0 18450
box 1578 1180 5350 3320
use bias_generator  bias_generator_12
timestamp 1722981971
transform 0 1 6220 -1 0 5850
box 1578 1180 5350 3320
use bias_generator  bias_generator_13
timestamp 1722981971
transform 0 1 6220 -1 0 10050
box 1578 1180 5350 3320
use bias_generator  bias_generator_14
timestamp 1722981971
transform 0 1 6220 -1 0 14250
box 1578 1180 5350 3320
use bias_generator  bias_generator_15
timestamp 1722981971
transform 0 1 6220 -1 0 18450
box 1578 1180 5350 3320
use sky130_fd_pr__pfet_01v8_8ND94H  sky130_fd_pr__pfet_01v8_8ND94H_0
timestamp 1722981971
transform 0 -1 3792 1 0 7723
box -123 -292 123 292
use sky130_fd_pr__pfet_01v8_8ND94H  sky130_fd_pr__pfet_01v8_8ND94H_1
timestamp 1722981971
transform 0 -1 3792 1 0 2523
box -123 -292 123 292
use sky130_fd_pr__pfet_01v8_8ND94H  sky130_fd_pr__pfet_01v8_8ND94H_2
timestamp 1722981971
transform 0 -1 3792 1 0 5123
box -123 -292 123 292
use sky130_fd_pr__pfet_01v8_8ND94H  sky130_fd_pr__pfet_01v8_8ND94H_3
timestamp 1722981971
transform 0 -1 3792 1 0 10323
box -123 -292 123 292
use sky130_fd_pr__pfet_01v8_8ND94H  sky130_fd_pr__pfet_01v8_8ND94H_4
timestamp 1722981971
transform 0 -1 3792 1 0 15523
box -123 -292 123 292
use sky130_fd_pr__pfet_01v8_8ND94H  sky130_fd_pr__pfet_01v8_8ND94H_5
timestamp 1722981971
transform 0 -1 3792 1 0 12923
box -123 -292 123 292
use sky130_fd_pr__pfet_01v8_8ND94H  sky130_fd_pr__pfet_01v8_8ND94H_6
timestamp 1722981971
transform 0 -1 3792 1 0 18123
box -123 -292 123 292
use sky130_fd_pr__pfet_01v8_8ND94H  sky130_fd_pr__pfet_01v8_8ND94H_7
timestamp 1722981971
transform 0 -1 3792 1 0 20723
box -123 -292 123 292
use sky130_fd_pr__pfet_01v8_8ND94H  sky130_fd_pr__pfet_01v8_8ND94H_8
timestamp 1722981971
transform 1 0 6823 0 1 1092
box -123 -292 123 292
use sky130_fd_pr__pfet_01v8_8ND94H  sky130_fd_pr__pfet_01v8_8ND94H_9
timestamp 1722981971
transform 1 0 6823 0 1 5292
box -123 -292 123 292
use sky130_fd_pr__pfet_01v8_8ND94H  sky130_fd_pr__pfet_01v8_8ND94H_10
timestamp 1722981971
transform 1 0 9423 0 1 1092
box -123 -292 123 292
use sky130_fd_pr__pfet_01v8_8ND94H  sky130_fd_pr__pfet_01v8_8ND94H_11
timestamp 1722981971
transform 1 0 9423 0 1 5292
box -123 -292 123 292
use sky130_fd_pr__pfet_01v8_8ND94H  sky130_fd_pr__pfet_01v8_8ND94H_12
timestamp 1722981971
transform 1 0 6823 0 1 9492
box -123 -292 123 292
use sky130_fd_pr__pfet_01v8_8ND94H  sky130_fd_pr__pfet_01v8_8ND94H_13
timestamp 1722981971
transform 1 0 6823 0 1 13692
box -123 -292 123 292
use sky130_fd_pr__pfet_01v8_8ND94H  sky130_fd_pr__pfet_01v8_8ND94H_14
timestamp 1722981971
transform 1 0 9423 0 1 9492
box -123 -292 123 292
use sky130_fd_pr__pfet_01v8_8ND94H  sky130_fd_pr__pfet_01v8_8ND94H_15
timestamp 1722981971
transform 1 0 9423 0 1 13692
box -123 -292 123 292
<< labels >>
flabel metal4 s 14383 22476 14413 22576 0 FreeSans 240 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 14659 22476 14689 22576 0 FreeSans 240 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 14107 22476 14137 22576 0 FreeSans 240 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 15181 0 15271 100 0 FreeSans 480 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 13249 0 13339 100 0 FreeSans 480 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 11317 0 11407 100 0 FreeSans 480 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 9385 0 9475 100 0 FreeSans 480 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 7453 0 7543 100 0 FreeSans 480 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 5521 0 5611 100 0 FreeSans 480 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 3589 0 3679 100 0 FreeSans 480 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 1657 0 1747 100 0 FreeSans 480 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 13831 22476 13861 22576 0 FreeSans 240 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 13555 22476 13585 22576 0 FreeSans 240 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 13279 22476 13309 22576 0 FreeSans 240 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 13003 22476 13033 22576 0 FreeSans 240 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 12727 22476 12757 22576 0 FreeSans 240 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 12451 22476 12481 22576 0 FreeSans 240 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 12175 22476 12205 22576 0 FreeSans 240 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 11899 22476 11929 22576 0 FreeSans 240 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 11623 22476 11653 22576 0 FreeSans 240 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 11347 22476 11377 22576 0 FreeSans 240 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 11071 22476 11101 22576 0 FreeSans 240 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 10795 22476 10825 22576 0 FreeSans 240 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 10519 22476 10549 22576 0 FreeSans 240 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 10243 22476 10273 22576 0 FreeSans 240 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 9967 22476 9997 22576 0 FreeSans 240 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 9691 22476 9721 22576 0 FreeSans 240 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 4999 22476 5029 22576 0 FreeSans 240 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 4723 22476 4753 22576 0 FreeSans 240 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4447 22476 4477 22576 0 FreeSans 240 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 4171 22476 4201 22576 0 FreeSans 240 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3895 22476 3925 22576 0 FreeSans 240 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 3619 22476 3649 22576 0 FreeSans 240 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3343 22476 3373 22576 0 FreeSans 240 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3067 22476 3097 22576 0 FreeSans 240 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 7207 22476 7237 22576 0 FreeSans 240 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 6931 22476 6961 22576 0 FreeSans 240 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 6655 22476 6685 22576 0 FreeSans 240 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 6379 22476 6409 22576 0 FreeSans 240 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 6103 22476 6133 22576 0 FreeSans 240 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 5827 22476 5857 22576 0 FreeSans 240 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 5551 22476 5581 22576 0 FreeSans 240 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 5275 22476 5305 22576 0 FreeSans 240 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 9415 22476 9445 22576 0 FreeSans 240 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 9139 22476 9169 22576 0 FreeSans 240 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 8863 22476 8893 22576 0 FreeSans 240 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 8587 22476 8617 22576 0 FreeSans 240 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 8311 22476 8341 22576 0 FreeSans 240 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 8035 22476 8065 22576 0 FreeSans 240 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 7759 22476 7789 22576 0 FreeSans 240 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 7483 22476 7513 22576 0 FreeSans 240 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 100 500 300 22076 1 FreeSans 200 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 400 500 600 22076 1 FreeSans 200 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 16100 22576
<< end >>
