magic
tech sky130A
magscale 1 2
timestamp 1722872344
<< error_p >>
rect -29 445 29 451
rect -29 411 -17 445
rect -29 405 29 411
<< nwell >>
rect -246 -584 246 584
<< pmos >>
rect -50 -436 50 364
<< pdiff >>
rect -108 352 -50 364
rect -108 -424 -96 352
rect -62 -424 -50 352
rect -108 -436 -50 -424
rect 50 352 108 364
rect 50 -424 62 352
rect 96 -424 108 352
rect 50 -436 108 -424
<< pdiffc >>
rect -96 -424 -62 352
rect 62 -424 96 352
<< nsubdiff >>
rect -210 514 210 548
rect -210 -514 -176 514
rect 176 451 210 514
rect 176 -514 210 -451
rect -210 -548 210 -514
<< nsubdiffcont >>
rect 176 -451 210 451
<< poly >>
rect -50 445 50 461
rect -50 411 -34 445
rect 34 411 50 445
rect -50 364 50 411
rect -50 -462 50 -436
<< polycont >>
rect -34 411 34 445
<< locali >>
rect -210 514 210 548
rect -210 -514 -176 514
rect 176 451 210 514
rect -50 411 -34 445
rect 34 411 50 445
rect -96 352 -62 368
rect -96 -440 -62 -424
rect 62 352 96 368
rect 62 -440 96 -424
rect 176 -514 210 -451
rect -210 -548 210 -514
<< viali >>
rect -17 411 17 445
rect -96 -424 -62 352
rect 62 -424 96 352
rect 176 -257 210 257
<< metal1 >>
rect -29 445 29 451
rect -29 411 -17 445
rect 17 411 29 445
rect -29 405 29 411
rect -102 352 -56 364
rect -102 -424 -96 352
rect -62 -424 -56 352
rect -102 -436 -56 -424
rect 56 352 102 364
rect 56 -424 62 352
rect 96 -424 102 352
rect 170 257 216 269
rect 170 -257 176 257
rect 210 -257 216 257
rect 170 -269 216 -257
rect 56 -436 102 -424
<< properties >>
string FIXED_BBOX -193 -531 193 531
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4.0 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 0 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 50 viagl 0 viagt 0
<< end >>
